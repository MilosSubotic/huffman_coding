...
architecture ...
	...
	
	signal state      : t_states;
	signal next_state : t_states;

	...
begin
	...