...
architecture ...

	type t_states is (
		NEW_CHAR,
		UPPER_NIBBLE,
		LAST_STAGE
	);
	
	...
	
begin
	...
	